library verilog;
use verilog.vl_types.all;
entity sub_13_0 is
    port(
        cin             : in     vl_logic;
        a               : in     vl_logic_vector(12 downto 0);
        b               : in     vl_logic_vector(12 downto 0);
        d               : out    vl_logic_vector(12 downto 0);
        cout            : out    vl_logic;
        \p_r15_0_\      : in     vl_logic
    );
end sub_13_0;
